--***************--\
-- <SHIFTER.VHD> -- 
--***************--/

entity Shifter is
--	port(
--		
--	);
end Shifter;



architecture Behavioral of Shifter is
begin

--process()
--begin
--	
--
--	
--end process;

end Behavioral;
