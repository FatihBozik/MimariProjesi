--***************----\
-- <CONSTANTS.VHD> -- 
--***************----/

package Constants is

--global
constant width : natural := 32;	
constant regfile_depth : positive := 32;
constant regfile_adrsize : positive := 5;

end Constants;
