--library ieee;
--use ieee.numeric_std.all;
--use work.Constants.all;
--use ieee.std_logic_1164.all;
--
--
--package Functions is
--
--procedure clearReg(r : in register_array);
--	
--end package Functions;
--
--
--
--package body Functions is
--
--procedure clearReg(r : in register_array) is
--begin
--	
--end clearReg;
--
--end package body Functions;